module game1_fsm(input logic clk, output logic led, output logic hex);

endmodule